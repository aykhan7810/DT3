///////////////////////////////////////////////////////////
//
// Class: apb_sequencer
//
///////////////////////////////////////////////////////////

typedef uvm_sequencer #(apb_transaction) apb_sequencer;

