///////////////////////////////////////////////////////////
//
// Class: apb_sequence_config
//
///////////////////////////////////////////////////////////

class apb_sequence_config extends uvm_object;
   int apb_test_cycles;
endclass 
