package control_unit_env_pkg;

`ifndef SYNTHESIS
   
`include "uvm_macros.svh"

   import uvm_pkg::*;
   import apb_pkg::*;
   import apb_env_pkg::*;

`include "irq_transaction.svh"
`include "irq_monitor.svh"
`include "irq_agent.svh"   
`include "control_unit_agent.svh"
`include "control_unit_env.svh"   
   
`endif //  `ifndef SYNTHESIS
   
endpackage

   
